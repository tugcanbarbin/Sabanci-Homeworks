`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   05:46:45 12/15/2020
// Design Name:   CLA
// Module Name:   C:/Xilinx/TugcanBarbin_25168_lab2/CLA/testttt2.v
// Project Name:  CLA
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: CLA
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module testttt2;

	// Inputs
	reg [19:0] A;
	reg [19:0] B;
	reg Cin;

	// Outputs
	wire Carry;
	wire [19:0] Sum;

	// Instantiate the Unit Under Test (UUT)
	CLA uut (
		.A(A), 
		.B(B), 
		.Cin(Cin), 
		.Carry(Carry), 
		.Sum(Sum)
	);

	initial begin
		// Initialize Inputs
		A = 0;
		B = 0;
		Cin = 0;

		// Wait 100 ns for global reset to finish
		#100;
        
		// Add stimulus here
		A[0] = 1;
		A[1] = 1;
		A[2] = 0;
		A[3] = 0;
		A[4] = 0;
		A[5] = 1;
		A[6] = 0;
		A[7] = 0;
		A[8] = 0;
		A[9] = 0;
		A[10] = 0;
		A[11] = 0;
		A[12] = 1;
		A[13] = 0;
		A[14] = 0;
		A[15] = 0;
		A[16] = 0;
		A[17] = 1;
		A[18] = 0;
		A[19] = 0;
		B[0] = 0;
		B[1] = 0;
		B[2] = 0;
		B[3] = 1;
		B[4] = 1;
		B[5] = 1;
		B[6] = 0;
		B[7] = 0;
		B[8] = 1;
		B[9] = 0;
		B[10] = 0;
		B[11] = 0;
		B[12] = 1;
		B[13] = 0;
		B[14] = 0;
		B[15] = 0;
		B[16] = 0;
		B[17] = 0;
		B[18] = 0;
		B[19] = 0;
		Cin=0;
		#100;
		A[0] = 1;
		A[1] = 1;
		A[2] = 1;
		A[3] = 0;
		A[4] = 0;
		A[5] = 1;
		A[6] = 0;
		A[7] = 0;
		A[8] = 0;
		A[9] = 0;
		A[10] = 1;
		A[11] = 1;
		A[12] = 1;
		A[13] = 0;
		A[14] = 0;
		A[15] = 0;
		A[16] = 0;
		A[17] = 0;
		A[18] = 0;
		A[19] = 0;
		B[0] = 1;
		B[1] = 1;
		B[2] = 0;
		B[3] = 0;
		B[4] = 0;
		B[5] = 0;
		B[6] = 1;
		B[7] = 0;
		B[8] = 0;
		B[9] = 0;
		B[10] = 0;
		B[11] = 0;
		B[12] = 0;
		B[13] = 0;
		B[14] = 0;
		B[15] = 0;
		B[16] = 0;
		B[17] = 0;
		B[18] = 0;
		B[19] = 0;
		Cin=1;
		#100;
		A[0] = 1;
		A[1] = 0;
		A[2] = 0;
		A[3] = 0;
		A[4] = 0;
		A[5] = 0;
		A[6] = 0;
		A[7] = 0;
		A[8] = 0;
		A[9] = 0;
		A[10] = 0;
		A[11] = 0;
		A[12] = 0;
		A[13] = 0;
		A[14] = 0;
		A[15] = 0;
		A[16] = 1;
		A[17] = 0;
		A[18] = 0;
		A[19] = 0;
		B[0] = 1;
		B[1] = 1;
		B[2] = 0;
		B[3] = 0;
		B[4] = 1;
		B[5] = 0;
		B[6] = 0;
		B[7] = 0;
		B[8] = 0;
		B[9] = 0;
		B[10] = 0;
		B[11] = 0;
		B[12] = 1;
		B[13] = 1;
		B[14] = 1;
		B[15] = 1;
		B[16] = 1;
		B[17] = 0;
		B[18] = 0;
		B[19] = 0;
		Cin=0;
		#100;
		A[0] = 1;
		A[1] = 1;
		A[2] = 1;
		A[3] = 0;
		A[4] = 0;
		A[5] = 1;
		A[6] = 0;
		A[7] = 0;
		A[8] = 0;
		A[9] = 0;
		A[10] = 1;
		A[11] = 1;
		A[12] = 1;
		A[13] = 0;
		A[14] = 0;
		A[15] = 0;
		A[16] = 0;
		A[17] = 0;
		A[18] = 0;
		A[19] = 0;
		B[0] = 1;
		B[1] = 1;
		B[2] = 0;
		B[3] = 0;
		B[4] = 0;
		B[5] = 0;
		B[6] = 1;
		B[7] = 0;
		B[8] = 0;
		B[9] = 0;
		B[10] = 0;
		B[11] = 0;
		B[12] = 0;
		B[13] = 1;
		B[14] = 0;
		B[15] = 0;
		B[16] = 0;
		B[17] = 0;
		B[18] = 1;
		B[19] = 0;
		Cin=1;
		#100;
		A[0] = 1;
		A[1] = 1;
		A[2] = 1;
		A[3] = 0;
		A[4] = 0;
		A[5] = 1;
		A[6] = 0;
		A[7] = 0;
		A[8] = 0;
		A[9] = 0;
		A[10] = 1;
		A[11] = 1;
		A[12] = 1;
		A[13] = 0;
		A[14] = 0;
		A[15] = 0;
		A[16] = 0;
		A[17] = 0;
		A[18] = 0;
		A[19] = 0;
		B[0] = 1;
		B[1] = 1;
		B[2] = 0;
		B[3] = 0;
		B[4] = 0;
		B[5] = 0;
		B[6] = 1;
		B[7] = 0;
		B[8] = 0;
		B[9] = 0;
		B[10] = 0;
		B[11] = 0;
		B[12] = 0;
		B[13] = 1;
		B[14] = 0;
		B[15] = 0;
		B[16] = 0;
		B[17] = 0;
		B[18] = 1;
		B[19] = 0;
		Cin=0;
		#100;
		A[0] = 0;
		A[1] = 0;
		A[2] = 0;
		A[3] = 0;
		A[4] = 0;
		A[5] = 0;
		A[6] = 0;
		A[7] = 0;
		A[8] = 0;
		A[9] = 0;
		A[10] = 0;
		A[11] = 0;
		A[12] = 0;
		A[13] = 0;
		A[14] = 0;
		A[15] = 0;
		A[16] = 0;
		A[17] = 0;
		A[18] = 0;
		A[19] = 1;
		B[0] = 1;
		B[1] = 1;
		B[2] = 1;
		B[3] = 1;
		B[4] = 1;
		B[5] = 1;
		B[6] = 1;
		B[7] = 1;
		B[8] = 1;
		B[9] = 1;
		B[10] = 1;
		B[11] = 1;
		B[12] = 1;
		B[13] = 1;
		B[14] = 1;
		B[15] = 1;
		B[16] = 1;
		B[17] = 1;
		B[18] = 1;
		B[19] = 1;
		Cin=0;

	end
      
endmodule

